../v2_extended_txns/addr_types.svh