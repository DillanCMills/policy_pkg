../v4_embedded_policies/policy_base.svh