../v3_extended_policies/policy_base.svh