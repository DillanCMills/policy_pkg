../v2_extended_txns/testbench.sv