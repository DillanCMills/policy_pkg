../v1_original_policies/policy_base.svh