../v3_extended_policies/addr_types.svh