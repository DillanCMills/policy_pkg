../v4_embedded_policies/addr_types.svh